`include "defines.v"

module if_id(
    input wire                   rst,
    input wire                   clk,
    input wire [`INST_ADDR_BUS]  if_pc,
    input wire [`INST_BUS]       if_instr,
    input wire                   exception,
    input wire                   inst_stall,
    input wire                   stall,
	input wire [`EXCEP_TYPE_BUS] if_exception_type,
		
	output reg [`EXCEP_TYPE_BUS] id_exception_type,
    output reg [`INST_ADDR_BUS]  id_pc,
    output reg [`INST_BUS]       id_instr
    );
    
    always @ (posedge clk) begin
        if (rst == `RST_ENABLE || exception == `EXCEPTION_ON) begin
            id_pc <= `ZEROWORD32;
            id_instr <= `ZEROWORD32;
            id_exception_type <= 6'h0;
        end else begin
            if (stall == `NOSTOP) begin
                if (inst_stall == 1'b1) begin
                    id_pc <= `ZEROWORD32;
                    id_instr <= `ZEROWORD32;
                    id_exception_type <= `ZEROWORD32;
                end else begin
                    id_pc <= if_pc;
                    id_instr <= if_instr;
                    id_exception_type <= if_exception_type;
                end 
            end
        end
    end
endmodule
